entity beginning1 is
end entity;


architecture inside of beginning1 is
begin 

     process is
	  begin
	  
	  report"i love red";
	  
	  wait;
	  end process;
	  
end architecture inside;	  

